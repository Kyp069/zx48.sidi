
module clockctrl (
	inclk,
	ena,
	outclk);	

	input		inclk;
	input		ena;
	output		outclk;
endmodule
